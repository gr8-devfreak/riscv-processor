
`ifndef FILE_INCL
    `include "processor_defines.sv"
`endif

module decode_jump_inst(
    input logic [31:0] instruction_code,
    output logic [4:0] rd,
    output logic [4:0] rs1,
    output logic [20:0] imm,
    output logic [1:0] jump_control
);

// Edit the code here begin ---------------------------------------------------
    logic [6:0]opcode;
    logic [2:0]funct3;

    assign opcode=instruction_code[6:0];
    assign rd = instruction_code[11:7];
    assign funct3=instruction_code[14:12];
    
    always_comb begin
        if(opcode==7'b1101111) begin
            jump_control=`JAL;
            rs1=5'b0;
            imm={instruction_code[31],instruction_code[19:12],instruction_code[20],instruction_code[30:21],1'b0};
        end
        else if(opcode==7'b1100111 && funct3==3'h0) begin 
            jump_control=`JALR;
            rs1=instruction_code[19:15];
            imm=instruction_code[31:20] ;
        end
        else  begin
            rs1 = 5'b0;
            imm=21'b0;
            jump_control=`JMP_NOP;
        end
    end
// Edit the code here end -----------------------------------------------------

/*
	Following section is necessary for dumping waveforms. This is needed for debug and simulations
*/

`ifndef SUBMODULE_DISABLE_WAVES
    initial begin
        $dumpfile("./sim_build/decode_jump_inst.vcd");
        $dumpvars(0, decode_jump_inst);
    end
`endif

endmodule
